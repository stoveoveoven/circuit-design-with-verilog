module controller(s, reset, w, opcode, op, nsel, out);
    input s, reset;
    input[2:0] opcode;
    input[1:0] op;
    output w;
    output[2:0] nsel;
    output[] out;



endmodule