//top level module for the RISC
module labt_top();

endmodule

//a register, parameter specifies how many bits is stored
module reg()

endmodule

//Standard multiplexer
module MUX();

endmodule

//Shifter units that shifts left or right depending on input
module shifter();

endmodule

//a register with load enable
module regLoad();

endmodule

//Arithmetic Logic unit, handles ADD/SUB
module ALU();

endmodule

